library verilog;
use verilog.vl_types.all;
entity Memory256_16bits_tb is
end Memory256_16bits_tb;
