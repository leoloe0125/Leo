library verilog;
use verilog.vl_types.all;
entity Instruction_Decoder_tb is
end Instruction_Decoder_tb;
