library verilog;
use verilog.vl_types.all;
entity Controller_tb is
end Controller_tb;
