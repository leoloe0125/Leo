library verilog;
use verilog.vl_types.all;
entity Mux8to1_16bits_tb is
end Mux8to1_16bits_tb;
