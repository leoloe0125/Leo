library verilog;
use verilog.vl_types.all;
entity ALU_16bits_tb is
end ALU_16bits_tb;
