library verilog;
use verilog.vl_types.all;
entity FA_16bits_tb is
end FA_16bits_tb;
