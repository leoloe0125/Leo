library verilog;
use verilog.vl_types.all;
entity RF8_16bits_tb is
end RF8_16bits_tb;
