library verilog;
use verilog.vl_types.all;
entity Decoder3to8_tb is
end Decoder3to8_tb;
