library verilog;
use verilog.vl_types.all;
entity DFF_16bits_tb is
end DFF_16bits_tb;
